C:\MC12\data\al\Nyquist.CIR Transient Analysis
* Converted From Micro Cap Source file to PSPICE
*
V1 INTERIOR_NONE1 0 SIN (0 1 10MEG 0 0 0)
RV1 4 INTERIOR_NONE1 0.001 ;added by V1
X91 1 2 AMP
+PARAMS: GAIN=0.97
X92 2 3 F
+PARAMS: FS={EXP(-S*0.6)/POW(1+S*1.2,6)}
X95 4 5 1 SUM
+PARAMS: KA=1 KB=1
X96 4 5 F
+PARAMS: FS={1/(S*6.2)}
*
*
.SUBCKT AMP PINA PINB
+PARAMS: GAIN=1
E1 PINB 0 PINA 0 {GAIN}
RE1 PINA 0 1G;added by E1
.ENDS AMP
*
*
.SUBCKT F PINA PINB
+PARAMS: FS={1/(S+1K)}
E1 PINB 0 LAPLACE {V(PINA,0)} = {{FS}}
RE1 PINA 0 1G;added by E1
.ENDS F
*
*
.SUBCKT SUM PINA PINB PINC
+PARAMS: KA=1 KB=1
E1 PINC 0 VALUE = {{KA}*V(PINA)+{KB}*V(PINB)}
.ENDS SUM
*
.OPTIONS ACCT LIST OPTS ABSTOL=1pA CHGTOL=.01pC
+ DEFL=100u DEFW=100u
+ DIGDRVF=2
+ DIGDRVZ=20K DIGERRDEFAULT=20
+ DIGERRLIMIT=0 DIGFREQ=10GHz
+ DIGINITSTATE=0
+ DIGIOLVL=2 DIGMNTYMX=2 DIGMNTYSCALE=0.4
+ DIGOVRDRV=3 DIGTYMXSCALE=1.6
+ GMIN=1p
+ ITL1=100 ITL2=50 ITL4=10 PIVREL=1m PIVTOL=.1p
+ RELTOL=1m TNOM=27
+ TRTOL=7 VNTOL=1u
+ WIDTH=80
*
.LIB "C:\MC12\library\NOM.LIB"
*
.TEMP 27
.TRAN 3 150 0 UIC
.PRINT TRAN V(2)
.PLOT TRAN V(2)
.PRINT TRAN V(7)
.PLOT TRAN V(7)
.PROBE
.END
;$SpiceType=PSPICE